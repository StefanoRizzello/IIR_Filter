library verilog;
use verilog.vl_types.all;
entity tb_iir is
end tb_iir;
